module imem (
	input [15:0] addr,
	output [31:0] data
);

	reg [15:0] mem_rom [15:0];

endmodule
