module rv32pipe3 (results);

	wire [31:0] instruction;
	wire [4:0] address;
	wire clock, writeEn;

endmodule
