module controller (inst, ctrl)
	input		[16:0] inst;
	output	[0:10] ctrl;
	
	

endmodule